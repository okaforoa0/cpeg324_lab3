//program counter file
