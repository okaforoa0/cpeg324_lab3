library ieee;
use ieee.std_logic_1164.all;
--use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity main_alu is
    Port ( 
        A       : in  STD_LOGIC_VECTOR(15 downto 0);
        B       : in  STD_LOGIC_VECTOR(15 downto 0);
        clk     : in  STD_LOGIC;
        control : in  STD_LOGIC_VECTOR(1 downto 0);
        result  : out STD_LOGIC_VECTOR(15 downto 0)
    );
end main_alu;

architecture Behavioral of main_alu is

    -- internal signal to hold adder result
    signal adder_result : STD_LOGIC_VECTOR(15 downto 0);

    -- instantiate custom 16-bit adder
    component adder16bit
        Port (
            A   : in  STD_LOGIC_VECTOR(15 downto 0);
            B   : in  STD_LOGIC_VECTOR(15 downto 0);
            S   : out STD_LOGIC_VECTOR(15 downto 0)
        );
    end component;

begin

    -- adder instantiation
    U1: adder16bit port map (
        A => A,
        B => B,
        S => adder_result
    );

    -- ALU operations
    process(clk)
    begin
        if rising_edge(clk) then
            case control is
                when "00" => -- ADD
                    result <= adder_result;

                when "01" => -- SWAP halves of A
                    result <= A(7 downto 0) & A(15 downto 8);

                when "10" => -- FORWARD A
                    result <= A;

                when "11" => -- COMPARE lower halves
                    if (A(7 downto 0) = B(7 downto 0)) then
                        result <= (others => '0');
                        result(0) <= '1'; -- set bit 0 to 1 if equal
                    else
                        result <= (others => '0'); -- otherwise all zeros
                    end if;

                when others =>
                    result <= (others => '0');
            end case;
        end if;
    end process;

end Behavioral;